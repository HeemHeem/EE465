module delay(
    input sym_clk_ena, sam_clk_ena,
    output [1:0] symb_a
    output [1:0] delay_reg [2:0]

);








endmodule
module upsampler(   input clk,
                    input wire signed [17:0] sig_in,
                    output reg signed [17:0] sig_out);

// counter for upsampler
reg [1:0] counter;




always @ (posedge clk)





endmodule